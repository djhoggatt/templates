// template.sv
// Description of component


// Test Module
module template();

    // I/O
  
    // Constants

    // Registers
  
    // Assignment Logic

    // Transitional Logic

endmodule