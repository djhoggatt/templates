// templateTestBench.sv
// Description of test


// Test Module
module testBench;

    // I/O
  
    // Instantiation
    template TEMPLATE();
  
    // Initial setup
    initial
    begin

    end

    // Test
    initial
    begin

    end
  
    // Tasks
    task templateTask;
    begin

    end

endmodule